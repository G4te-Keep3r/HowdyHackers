LEF " Howdy Hackers "