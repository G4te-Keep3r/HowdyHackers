CkT " Howdy Hackers "