cDL " Howdy Hackers "