CdL " Howdy Hackers "