CKT " Howdy Hackers "