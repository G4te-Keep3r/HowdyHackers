lEF " Howdy Hackers "