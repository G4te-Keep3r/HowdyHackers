bsV " Howdy Hackers "