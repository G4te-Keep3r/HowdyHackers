VH " Howdy Hackers "