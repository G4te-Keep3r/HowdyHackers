sVH " Howdy Hackers "