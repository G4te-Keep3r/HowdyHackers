bSV " Howdy Hackers "