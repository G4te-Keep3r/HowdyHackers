vHD " Howdy Hackers "