BSV " Howdy Hackers "