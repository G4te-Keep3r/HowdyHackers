SV " Howdy Hackers "