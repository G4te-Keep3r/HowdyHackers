leF " Howdy Hackers "