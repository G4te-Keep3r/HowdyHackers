CDL " Howdy Hackers "