svH " Howdy Hackers "