cKT " Howdy Hackers "